`include "pkg.sv"
`include "tracer_pkg.sv"
`include "Program_Counter.sv"
`include "inst_mem.sv"
`include "mux_2x1.sv"
`include "mux_4x1.sv"
`include "pipe_reg.sv"
`include "hazard_detection.sv"
`include "Reg_file.sv"
`include "imm_gen.sv"
`include "Control_Unit.sv"
`include "Barrel_Shifter.sv"
`include "Flush.sv"
`include "branch_comp.sv"
`include "Branch_Selector.sv"
`include "alu_logic.sv"
`include "fwd_logic.sv"
`include "DMEM.sv"
`include "tracer.sv"
`include "Top.sv"